-- VHDL Test Fixture: Chain shift scenario
-- 8 registers at 0x00-0x1C for chain shift testing

library ieee;
use ieee.std_logic_1164.all;

entity addr_test_chain is
    port (
        clk : in std_logic;
        -- @axion BASE_ADDR=0x0000
        -- @axion RW ADDR=0x00
        chain_reg_0 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x04
        chain_reg_1 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x08
        chain_reg_2 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x0C
        chain_reg_3 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x10
        chain_reg_4 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x14
        chain_reg_5 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x18
        chain_reg_6 : inout std_logic_vector(31 downto 0);
        -- @axion RW ADDR=0x1C
        chain_reg_7 : inout std_logic_vector(31 downto 0)
    );
end entity addr_test_chain;

architecture rtl of addr_test_chain is
begin
end architecture rtl;
